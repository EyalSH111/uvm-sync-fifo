`include "fifo_if.sv"
`include "fifo_item.sv"



`include "fifo_driver.sv"
`include "fifo_monitor.sv"
`include "fifo_scoreboard.sv"
`include "fifo_coverage.sv"
`include "fifo_env.sv"

`include "fifo_random_test.sv"
`include "top_tb.sv"
`include "fifo_assertions.sv"
`include "fifo_reset_mid_test.sv"
